module controller(input logic ph1, ph2, reset,
                  output logic dataClk1, dataClk2, clearAccum,
                  output logic[1:0] muxControl );
endmodule