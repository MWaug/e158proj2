module controller(input logic clk1, clk2, reset,
                  output logic dataClk1, dataClk2, clearAccum,
                  output logic[1:0] muxControl );
endmodule